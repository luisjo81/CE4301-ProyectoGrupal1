module procesador()




endmodule
