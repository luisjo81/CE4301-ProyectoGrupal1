module tb_decoInst();

logic [25:0] inst;
clk = 0;

decoInst decoInst (.)

initial
begin



end


endmodule 