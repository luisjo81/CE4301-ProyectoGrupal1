module decoInst (input logic inst, output logic opcode);
$display("Mariano")




endmodule